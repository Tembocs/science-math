module main
// import math
import mathematics as mts

fn main() {
	fraction1 := mts.Fraction {
		8,
		7
	}

	println('Numerator: $fraction1.numerator')
	println('Numerator: $fraction1.denominator')
}