module main

import mathematics as mts

fn main() {
	some_numbers := [24, 36, 72]

	println('GCF of $some_numbers = ${mts.gcf(some_numbers)}')
}