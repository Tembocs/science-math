module main

import mathematics as mts

fn main() {
	some_numbers := [56, 112,210]
	println('Hello World!')
	println('The GCF of $some_numbers is ${mts.gcf(some_numbers)}')
}